module asc16x8 (
   input  wire        clk,
   input  wire [10:0]  bitmap_addr,
   output wire  [7:0]  bitmap_byte 
);


`ifdef SIM 
   reg [7:0]   bitmap_reg [ 0 : 2047 ] ; 
   reg         bitmap_byte_r ; 

   assign   bitmap_byte =  bitmap_byte_r ;   
   initial begin 
      $readmemh("../rtl/asc16x8.mem", bitmap_reg, 0, 2047 ) ;    
   end 

   always @( posedge clk ) begin  
      bitmap_byte_r <= bitmap_reg[ bitmap_addr] ;  
   end 
`else 
   
   asc16X8_xilinx asc16X8_xilinx_inst (
     .clka     (  clk         ), // input clka
     .addra    (  bitmap_addr ), // input [10 : 0] addra
     .douta    (  bitmap_byte )  // output [7 : 0] douta
   );


`endif 



endmodule   
/*******************************************************************************
*     This file is owned and controlled by Xilinx and must be used solely      *
*     for design, simulation, implementation and creation of design files      *
*     limited to Xilinx devices or technologies. Use with non-Xilinx           *
*     devices or technologies is expressly prohibited and immediately          *
*     terminates your license.                                                 *
*                                                                              *
*     XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY     *
*     FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY     *
*     PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE              *
*     IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS       *
*     MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY       *
*     CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY        *
*     RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY        *
*     DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE    *
*     IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR           *
*     REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF          *
*     INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A    *
*     PARTICULAR PURPOSE.                                                      *
*                                                                              *
*     Xilinx products are not intended for use in life support appliances,     *
*     devices, or systems.  Use in such applications are expressly             *
*     prohibited.                                                              *
*                                                                              *
*     (c) Copyright 1995-2014 Xilinx, Inc.                                     *
*     All rights reserved.                                                     *
*******************************************************************************/

/*******************************************************************************
*     Generated from core with identifier: xilinx.com:ip:blk_mem_gen:7.3       *
*                                                                              *
*     The Xilinx LogiCORE IP Block Memory Generator replaces the Dual Port     *
*     Block Memory and Single Port Block Memory LogiCOREs, but is not a        *
*     direct drop-in replacement.  It should be used in all new Xilinx         *
*     designs. The core supports RAM and ROM functions over a wide range of    *
*     widths and depths. Use this core to generate block memories with         *
*     symmetric or asymmetric read and write port widths, as well as cores     *
*     which can perform simultaneous write operations to separate              *
*     locations, and simultaneous read operations from the same location.      *
*     For more information on differences in interface and feature support     *
*     between this core and the Dual Port Block Memory and Single Port         *
*     Block Memory LogiCOREs, please consult the data sheet.                   *
*******************************************************************************/

// The following must be inserted into your Verilog file for this
// core to be instantiated. Change the instance name and port connections
// (in parentheses) to your own signal names.

//----------- Begin Cut here for INSTANTIATION Template ---// INST_TAG
// INST_TAG_END ------ End INSTANTIATION Template ---------

// You must compile the wrapper file asc16X8_xilinx.v when simulating
// the core, asc16X8_xilinx. When compiling the wrapper file, be sure to
// reference the XilinxCoreLib Verilog simulation library. For detailed
// instructions, please refer to the "CORE Generator Help".

