
parameter BLACK = 3'b000; 
parameter BLUE  = 3'b001; 
parameter GREEN = 3'b010; 
parameter CYAN  = 3'b011; 
parameter RED   = 3'b100; 
parameter MAGENTA  = 3'b101; 
parameter YELLOW = 3'b110; 
parameter WHITE = 3'b111; 


parameter TEXT_LOGO_BIT  = 0; 
parameter TEXT_SCORE_BIT = 1; 
parameter TEXT_OVER_BIT  = 2; 
